// Decoder for


module corrector (input [271:0] IN,
    input [15:0] SYN,
    output logic [271:0] OUT
);

logic [271:0] LOC;

    always_comb begin
       case (SYN)
        16'b0100111100001001 : LOC = 272'd1 << 0 ;
        16'b1110011101000110 : LOC = 272'd1 << 1 ;
        16'b0101010111111000 : LOC = 272'd1 << 2 ;
        16'b0011001001110100 : LOC = 272'd1 << 3 ;
        16'b0111100000011001 : LOC = 272'd1 << 4 ;
        16'b0010010010010111 : LOC = 272'd1 << 5 ;
        16'b0010110111011001 : LOC = 272'd1 << 6 ;
        16'b1010000110100011 : LOC = 272'd1 << 7 ;
        16'b0000011011110001 : LOC = 272'd1 << 8 ;
        16'b0001011101011110 : LOC = 272'd1 << 9 ;
        16'b0000110111001100 : LOC = 272'd1 << 10 ;
        16'b1001110001011011 : LOC = 272'd1 << 11 ;
        16'b1101010110010000 : LOC = 272'd1 << 12 ;
        16'b1010001000111001 : LOC = 272'd1 << 13 ;
        16'b0010010010101101 : LOC = 272'd1 << 14 ;
        16'b1101101011101000 : LOC = 272'd1 << 15 ;
        16'b0000010000011101 : LOC = 272'd1 << 16 ;
        16'b0010111100100010 : LOC = 272'd1 << 17 ;
        16'b1011000010000111 : LOC = 272'd1 << 18 ;
        16'b0001111011011010 : LOC = 272'd1 << 19 ;
        16'b1111000101100000 : LOC = 272'd1 << 20 ;
        16'b0000100101011011 : LOC = 272'd1 << 21 ;
        16'b0000110011010000 : LOC = 272'd1 << 22 ;
        16'b1011011010010110 : LOC = 272'd1 << 23 ;
        16'b1010011111110000 : LOC = 272'd1 << 24 ;
        16'b1100010100101001 : LOC = 272'd1 << 25 ;
        16'b1000101110001001 : LOC = 272'd1 << 26 ;
        16'b0000110110110111 : LOC = 272'd1 << 27 ;
        16'b0001111011101001 : LOC = 272'd1 << 28 ;
        16'b0111010001011000 : LOC = 272'd1 << 29 ;
        16'b0010101101110110 : LOC = 272'd1 << 30 ;
        16'b0010111010100111 : LOC = 272'd1 << 31 ;
        16'b1101101000011011 : LOC = 272'd1 << 32 ;
        16'b0110011000000001 : LOC = 272'd1 << 33 ;
        16'b0000111010011001 : LOC = 272'd1 << 34 ;
        16'b1111110010101000 : LOC = 272'd1 << 35 ;
        16'b1000110000100001 : LOC = 272'd1 << 36 ;
        16'b0100100011101001 : LOC = 272'd1 << 37 ;
        16'b1100000111100111 : LOC = 272'd1 << 38 ;
        16'b1011001101110111 : LOC = 272'd1 << 39 ;
        16'b1011100000100011 : LOC = 272'd1 << 40 ;
        16'b0110101001010100 : LOC = 272'd1 << 41 ;
        16'b1000001101011100 : LOC = 272'd1 << 42 ;
        16'b0101100001010110 : LOC = 272'd1 << 43 ;
        16'b1100101011010011 : LOC = 272'd1 << 44 ;
        16'b0011111100001011 : LOC = 272'd1 << 45 ;
        16'b0001010011001110 : LOC = 272'd1 << 46 ;
        16'b1000010110111011 : LOC = 272'd1 << 47 ;
        16'b1101001110011100 : LOC = 272'd1 << 48 ;
        16'b0010011100001000 : LOC = 272'd1 << 49 ;
        16'b1111110000000100 : LOC = 272'd1 << 50 ;
        16'b1100111100010101 : LOC = 272'd1 << 51 ;
        16'b1011100100100100 : LOC = 272'd1 << 52 ;
        16'b0111101011110110 : LOC = 272'd1 << 53 ;
        16'b1001101001010100 : LOC = 272'd1 << 54 ;
        16'b0110010101101101 : LOC = 272'd1 << 55 ;
        16'b0101100101111100 : LOC = 272'd1 << 56 ;
        16'b0000110000100110 : LOC = 272'd1 << 57 ;
        16'b1011111011000010 : LOC = 272'd1 << 58 ;
        16'b0110010011000011 : LOC = 272'd1 << 59 ;
        16'b0000011001010111 : LOC = 272'd1 << 60 ;
        16'b0111001101110001 : LOC = 272'd1 << 61 ;
        16'b1001011100010010 : LOC = 272'd1 << 62 ;
        16'b0001000101101110 : LOC = 272'd1 << 63 ;
        16'b0110000110010011 : LOC = 272'd1 << 64 ;
        16'b0001111110000010 : LOC = 272'd1 << 65 ;
        16'b0001001000010101 : LOC = 272'd1 << 66 ;
        16'b1110111010000000 : LOC = 272'd1 << 67 ;
        16'b1110010000010000 : LOC = 272'd1 << 68 ;
        16'b0111001100101011 : LOC = 272'd1 << 69 ;
        16'b1001010111010101 : LOC = 272'd1 << 70 ;
        16'b1010011101101100 : LOC = 272'd1 << 71 ;
        16'b1010010010000001 : LOC = 272'd1 << 72 ;
        16'b0101100100010011 : LOC = 272'd1 << 73 ;
        16'b1000001110110010 : LOC = 272'd1 << 74 ;
        16'b0011100110100001 : LOC = 272'd1 << 75 ;
        16'b1011100011000100 : LOC = 272'd1 << 76 ;
        16'b0101100010100101 : LOC = 272'd1 << 77 ;
        16'b1000111011001110 : LOC = 272'd1 << 78 ;
        16'b1100101010100100 : LOC = 272'd1 << 79 ;
        16'b1010100000001010 : LOC = 272'd1 << 80 ;
        16'b0001001100001001 : LOC = 272'd1 << 81 ;
        16'b1011011011011000 : LOC = 272'd1 << 82 ;
        16'b0110011111011011 : LOC = 272'd1 << 83 ;
        16'b0101110101010000 : LOC = 272'd1 << 84 ;
        16'b1011000001001101 : LOC = 272'd1 << 85 ;
        16'b1011010000011010 : LOC = 272'd1 << 86 ;
        16'b0100110001001011 : LOC = 272'd1 << 87 ;
        16'b1110000011101101 : LOC = 272'd1 << 88 ;
        16'b0010000101100010 : LOC = 272'd1 << 89 ;
        16'b0001100011110100 : LOC = 272'd1 << 90 ;
        16'b1110001011010000 : LOC = 272'd1 << 91 ;
        16'b1000111010000101 : LOC = 272'd1 << 92 ;
        16'b0101010010010110 : LOC = 272'd1 << 93 ;
        16'b0110110011010110 : LOC = 272'd1 << 94 ;
        16'b0011000100111010 : LOC = 272'd1 << 95 ;
        16'b0001000111001011 : LOC = 272'd1 << 96 ;
        16'b1011000111000001 : LOC = 272'd1 << 97 ;
        16'b0111101001100000 : LOC = 272'd1 << 98 ;
        16'b1000111010101000 : LOC = 272'd1 << 99 ;
        16'b0100010100110000 : LOC = 272'd1 << 100 ;
        16'b1001101111000110 : LOC = 272'd1 << 101 ;
        16'b1101000000001001 : LOC = 272'd1 << 102 ;
        16'b0101011110110001 : LOC = 272'd1 << 103 ;
        16'b1101000101000110 : LOC = 272'd1 << 104 ;
        16'b1100110110000100 : LOC = 272'd1 << 105 ;
        16'b0100111011100011 : LOC = 272'd1 << 106 ;
        16'b0010011110100001 : LOC = 272'd1 << 107 ;
        16'b0001110011011101 : LOC = 272'd1 << 108 ;
        16'b0011000100010001 : LOC = 272'd1 << 109 ;
        16'b1010010011001100 : LOC = 272'd1 << 110 ;
        16'b1101100110011010 : LOC = 272'd1 << 111 ;
        16'b1010011110000010 : LOC = 272'd1 << 112 ;
        16'b1000100000111011 : LOC = 272'd1 << 113 ;
        16'b0110100101001001 : LOC = 272'd1 << 114 ;
        16'b0110101010001001 : LOC = 272'd1 << 115 ;
        16'b0101011101011001 : LOC = 272'd1 << 116 ;
        16'b0100110010001110 : LOC = 272'd1 << 117 ;
        16'b1100011001101000 : LOC = 272'd1 << 118 ;
        16'b0011010011100010 : LOC = 272'd1 << 119 ;
        16'b0011010110000000 : LOC = 272'd1 << 120 ;
        16'b0010001101010101 : LOC = 272'd1 << 121 ;
        16'b0011100010010101 : LOC = 272'd1 << 122 ;
        16'b0010000001011010 : LOC = 272'd1 << 123 ;
        16'b0000000011100011 : LOC = 272'd1 << 124 ;
        16'b0100001100010010 : LOC = 272'd1 << 125 ;
        16'b0110100010110010 : LOC = 272'd1 << 126 ;
        16'b0001010001100111 : LOC = 272'd1 << 127 ;
        16'b1000101110100111 : LOC = 272'd1 << 128 ;
        16'b1100110011000001 : LOC = 272'd1 << 129 ;
        16'b1100010001110001 : LOC = 272'd1 << 130 ;
        16'b1011000001111011 : LOC = 272'd1 << 131 ;
        16'b0001110000010010 : LOC = 272'd1 << 132 ;
        16'b0100011001001101 : LOC = 272'd1 << 133 ;
        16'b0000000011011100 : LOC = 272'd1 << 134 ;
        16'b0011100101000011 : LOC = 272'd1 << 135 ;
        16'b1000001010000011 : LOC = 272'd1 << 136 ;
        16'b1001000000010110 : LOC = 272'd1 << 137 ;
        16'b1001000100000101 : LOC = 272'd1 << 138 ;
        16'b0001001010110110 : LOC = 272'd1 << 139 ;
        16'b0000100001110001 : LOC = 272'd1 << 140 ;
        16'b0110000110100000 : LOC = 272'd1 << 141 ;
        16'b1011011000000000 : LOC = 272'd1 << 142 ;
        16'b1011111001001100 : LOC = 272'd1 << 143 ;
        16'b0100001010000101 : LOC = 272'd1 << 144 ;
        16'b0110010111000100 : LOC = 272'd1 << 145 ;
        16'b0000010101001111 : LOC = 272'd1 << 146 ;
        16'b1000000001110111 : LOC = 272'd1 << 147 ;
        16'b1100000100100100 : LOC = 272'd1 << 148 ;
        16'b0001001101010000 : LOC = 272'd1 << 149 ;
        16'b1011001011100000 : LOC = 272'd1 << 150 ;
        16'b1110100111100010 : LOC = 272'd1 << 151 ;
        16'b0010100000011100 : LOC = 272'd1 << 152 ;
        16'b0100000000111001 : LOC = 272'd1 << 153 ;
        16'b0010001010101011 : LOC = 272'd1 << 154 ;
        16'b1110111100011000 : LOC = 272'd1 << 155 ;
        16'b0001000000001111 : LOC = 272'd1 << 156 ;
        16'b0000111101011000 : LOC = 272'd1 << 157 ;
        16'b0011100000101101 : LOC = 272'd1 << 158 ;
        16'b0100001101100101 : LOC = 272'd1 << 159 ;
        16'b0101001000001100 : LOC = 272'd1 << 160 ;
        16'b0101101010101110 : LOC = 272'd1 << 161 ;
        16'b0100000111110010 : LOC = 272'd1 << 162 ;
        16'b0100101000111100 : LOC = 272'd1 << 163 ;
        16'b1100010010011001 : LOC = 272'd1 << 164 ;
        16'b1111000110000100 : LOC = 272'd1 << 165 ;
        16'b0000010001111000 : LOC = 272'd1 << 166 ;
        16'b0000100010000111 : LOC = 272'd1 << 167 ;
        16'b1001000100111100 : LOC = 272'd1 << 168 ;
        16'b0001010100010100 : LOC = 272'd1 << 169 ;
        16'b0001100110101100 : LOC = 272'd1 << 170 ;
        16'b0101100010000010 : LOC = 272'd1 << 171 ;
        16'b0110100100101010 : LOC = 272'd1 << 172 ;
        16'b0001101010001000 : LOC = 272'd1 << 173 ;
        16'b0010010100000110 : LOC = 272'd1 << 174 ;
        16'b0010000001101001 : LOC = 272'd1 << 175 ;
        16'b0101010000100100 : LOC = 272'd1 << 176 ;
        16'b0010010001010001 : LOC = 272'd1 << 177 ;
        16'b1100001000011000 : LOC = 272'd1 << 178 ;
        16'b0001100100001010 : LOC = 272'd1 << 179 ;
        16'b1100111000001100 : LOC = 272'd1 << 180 ;
        16'b0000000111000101 : LOC = 272'd1 << 181 ;
        16'b0111111000001000 : LOC = 272'd1 << 182 ;
        16'b1001110000101100 : LOC = 272'd1 << 183 ;
        16'b1001010000100010 : LOC = 272'd1 << 184 ;
        16'b1010000011000010 : LOC = 272'd1 << 185 ;
        16'b0100000100101111 : LOC = 272'd1 << 186 ;
        16'b0010001010010001 : LOC = 272'd1 << 187 ;
        16'b1001000011010000 : LOC = 272'd1 << 188 ;
        16'b0101011000110111 : LOC = 272'd1 << 189 ;
        16'b1100000010001100 : LOC = 272'd1 << 190 ;
        16'b0100000001110100 : LOC = 272'd1 << 191 ;
        16'b1111100001000010 : LOC = 272'd1 << 192 ;
        16'b0100111011000100 : LOC = 272'd1 << 193 ;
        16'b0000010010001011 : LOC = 272'd1 << 194 ;
        16'b0011001000101110 : LOC = 272'd1 << 195 ;
        16'b0111000011000000 : LOC = 272'd1 << 196 ;
        16'b0100011001000010 : LOC = 272'd1 << 197 ;
        16'b0110001100000100 : LOC = 272'd1 << 198 ;
        16'b0011100000000110 : LOC = 272'd1 << 199 ;
        16'b0001011001000001 : LOC = 272'd1 << 200 ;
        16'b0100000100011100 : LOC = 272'd1 << 201 ;
        16'b0000100100010101 : LOC = 272'd1 << 202 ;
        16'b1000100100000110 : LOC = 272'd1 << 203 ;
        16'b0010110001000010 : LOC = 272'd1 << 204 ;
        16'b0000011000100011 : LOC = 272'd1 << 205 ;
        16'b0101110010011000 : LOC = 272'd1 << 206 ;
        16'b0110011101100000 : LOC = 272'd1 << 207 ;
        16'b0101100100000100 : LOC = 272'd1 << 208 ;
        16'b0010101010000010 : LOC = 272'd1 << 209 ;
        16'b1000101010011100 : LOC = 272'd1 << 210 ;
        16'b0100000101010001 : LOC = 272'd1 << 211 ;
        16'b0101101011000001 : LOC = 272'd1 << 212 ;
        16'b1100100110101000 : LOC = 272'd1 << 213 ;
        16'b0011101000010000 : LOC = 272'd1 << 214 ;
        16'b1000101111100000 : LOC = 272'd1 << 215 ;
        16'b0000101000010110 : LOC = 272'd1 << 216 ;
        16'b1101000001100101 : LOC = 272'd1 << 217 ;
        16'b1000000010110100 : LOC = 272'd1 << 218 ;
        16'b0100100111000000 : LOC = 272'd1 << 219 ;
        16'b1000010000010011 : LOC = 272'd1 << 220 ;
        16'b0001100101100000 : LOC = 272'd1 << 221 ;
        16'b0011010000001001 : LOC = 272'd1 << 222 ;
        16'b1110000100000010 : LOC = 272'd1 << 223 ;
        16'b1000010110100000 : LOC = 272'd1 << 224 ;
        16'b0101001000100001 : LOC = 272'd1 << 225 ;
        16'b0100001010101000 : LOC = 272'd1 << 226 ;
        16'b0100101000001010 : LOC = 272'd1 << 227 ;
        16'b0000011001100100 : LOC = 272'd1 << 228 ;
        16'b0000011011001000 : LOC = 272'd1 << 229 ;
        16'b0101000001101000 : LOC = 272'd1 << 230 ;
        16'b1101100011011001 : LOC = 272'd1 << 231 ;
        16'b0011000101001000 : LOC = 272'd1 << 232 ;
        16'b0101101110010000 : LOC = 272'd1 << 233 ;
        16'b0110000010110101 : LOC = 272'd1 << 234 ;
        16'b0000000110010110 : LOC = 272'd1 << 235 ;
        16'b1001000001000011 : LOC = 272'd1 << 236 ;
        16'b0010011000010010 : LOC = 272'd1 << 237 ;
        16'b0000001110100100 : LOC = 272'd1 << 238 ;
        16'b1010001100010000 : LOC = 272'd1 << 239 ;
        16'b0001000110011000 : LOC = 272'd1 << 240 ;
        16'b1000100000001101 : LOC = 272'd1 << 241 ;
        16'b0001100001001001 : LOC = 272'd1 << 242 ;
        16'b0001000010110001 : LOC = 272'd1 << 243 ;
        16'b0010000000100111 : LOC = 272'd1 << 244 ;
        16'b0000010100100101 : LOC = 272'd1 << 245 ;
        16'b1100000010100010 : LOC = 272'd1 << 246 ;
        16'b1010100010100000 : LOC = 272'd1 << 247 ;
        16'b0001000010101010 : LOC = 272'd1 << 248 ;
        16'b0000001000101101 : LOC = 272'd1 << 249 ;
        16'b1000111100000000 : LOC = 272'd1 << 250 ;
        16'b0110010000101000 : LOC = 272'd1 << 251 ;
        16'b0100000001001110 : LOC = 272'd1 << 252 ;
        16'b1100000000010101 : LOC = 272'd1 << 253 ;
        16'b1010101000000100 : LOC = 272'd1 << 254 ;
        16'b0001110010100000 : LOC = 272'd1 << 255 ;
        16'b0000000000000001 : LOC = 272'd1 << 256 ;
        16'b0000000000000010 : LOC = 272'd1 << 257 ;
        16'b0000000000000100 : LOC = 272'd1 << 258 ;
        16'b0000000000001000 : LOC = 272'd1 << 259 ;
        16'b0000000000010000 : LOC = 272'd1 << 260 ;
        16'b0000000000100000 : LOC = 272'd1 << 261 ;
        16'b0000000001000000 : LOC = 272'd1 << 262 ;
        16'b0000000010000000 : LOC = 272'd1 << 263 ;
        16'b0000000100000000 : LOC = 272'd1 << 264 ;
        16'b0000001000000000 : LOC = 272'd1 << 265 ;
        16'b0000010000000000 : LOC = 272'd1 << 266 ;
        16'b0000100000000000 : LOC = 272'd1 << 267 ;
        16'b0001000000000000 : LOC = 272'd1 << 268 ;
        16'b0010000000000000 : LOC = 272'd1 << 269 ;
        16'b0100000000000000 : LOC = 272'd1 << 270 ;
        16'b1000000000000000 : LOC = 272'd1 << 271 ;
        default: LOC = 272'd0;
        endcase
        OUT = IN ^ LOC ;
    end
endmodule


module dec_top (
    input [271:0] IN,
    output wire [271:0] OUT,
    output reg [15:0] SYN,
    output reg ERR, SGL, DBL
);

    wire [15:0] CHK = IN[271:256];

    always_comb begin
        SYN[0] = IN[0] ^ IN[4] ^ IN[5] ^ IN[6] ^ IN[7] ^ IN[8] ^ IN[11] ^ IN[13] ^ IN[14] ^ IN[16] ^ IN[18] ^ IN[21] ^ IN[25] ^ IN[26] ^ IN[27] ^ IN[28] ^ IN[31] ^ IN[32] ^ IN[33] ^ IN[34] ^ IN[36] ^ IN[37] ^ IN[38] ^ IN[39] ^ IN[40] ^ IN[44] ^ IN[45] ^ IN[47] ^ IN[51] ^ IN[55] ^ IN[59] ^ IN[60] ^ IN[61] ^ IN[64] ^ IN[66] ^ IN[69] ^ IN[70] ^ IN[72] ^ IN[73] ^ IN[75] ^ IN[77] ^ IN[81] ^ IN[83] ^ IN[85] ^ IN[87] ^ IN[88] ^ IN[92] ^ IN[96] ^ IN[97] ^ IN[102] ^ IN[103] ^ IN[106] ^ IN[107] ^ IN[108] ^ IN[109] ^ IN[113] ^ IN[114] ^ IN[115] ^ IN[116] ^ IN[121] ^ IN[122] ^ IN[124] ^ IN[127] ^ IN[128] ^ IN[129] ^ IN[130] ^ IN[131] ^ IN[133] ^ IN[135] ^ IN[136] ^ IN[138] ^ IN[140] ^ IN[144] ^ IN[146] ^ IN[147] ^ IN[153] ^ IN[154] ^ IN[156] ^ IN[158] ^ IN[159] ^ IN[164] ^ IN[167] ^ IN[175] ^ IN[177] ^ IN[181] ^ IN[186] ^ IN[187] ^ IN[189] ^ IN[194] ^ IN[200] ^ IN[202] ^ IN[205] ^ IN[211] ^ IN[212] ^ IN[217] ^ IN[220] ^ IN[222] ^ IN[225] ^ IN[231] ^ IN[234] ^ IN[236] ^ IN[241] ^ IN[242] ^ IN[243] ^ IN[244] ^ IN[245] ^ IN[249] ^ IN[253] ^ CHK[0];
        SYN[1] = IN[1] ^ IN[5] ^ IN[7] ^ IN[9] ^ IN[11] ^ IN[17] ^ IN[18] ^ IN[19] ^ IN[21] ^ IN[23] ^ IN[27] ^ IN[30] ^ IN[31] ^ IN[32] ^ IN[38] ^ IN[39] ^ IN[40] ^ IN[43] ^ IN[44] ^ IN[45] ^ IN[46] ^ IN[47] ^ IN[53] ^ IN[57] ^ IN[58] ^ IN[59] ^ IN[60] ^ IN[62] ^ IN[63] ^ IN[64] ^ IN[65] ^ IN[69] ^ IN[73] ^ IN[74] ^ IN[78] ^ IN[80] ^ IN[83] ^ IN[86] ^ IN[87] ^ IN[89] ^ IN[93] ^ IN[94] ^ IN[95] ^ IN[96] ^ IN[101] ^ IN[104] ^ IN[106] ^ IN[111] ^ IN[112] ^ IN[113] ^ IN[117] ^ IN[119] ^ IN[123] ^ IN[124] ^ IN[125] ^ IN[126] ^ IN[127] ^ IN[128] ^ IN[131] ^ IN[132] ^ IN[135] ^ IN[136] ^ IN[137] ^ IN[139] ^ IN[146] ^ IN[147] ^ IN[151] ^ IN[154] ^ IN[156] ^ IN[161] ^ IN[162] ^ IN[167] ^ IN[171] ^ IN[172] ^ IN[174] ^ IN[179] ^ IN[184] ^ IN[185] ^ IN[186] ^ IN[189] ^ IN[192] ^ IN[194] ^ IN[195] ^ IN[197] ^ IN[199] ^ IN[203] ^ IN[204] ^ IN[205] ^ IN[209] ^ IN[216] ^ IN[220] ^ IN[223] ^ IN[227] ^ IN[235] ^ IN[236] ^ IN[237] ^ IN[244] ^ IN[246] ^ IN[248] ^ IN[252] ^ CHK[1];
        SYN[2] = IN[1] ^ IN[3] ^ IN[5] ^ IN[9] ^ IN[10] ^ IN[14] ^ IN[16] ^ IN[18] ^ IN[23] ^ IN[27] ^ IN[30] ^ IN[31] ^ IN[38] ^ IN[39] ^ IN[41] ^ IN[42] ^ IN[43] ^ IN[46] ^ IN[48] ^ IN[50] ^ IN[51] ^ IN[52] ^ IN[53] ^ IN[54] ^ IN[55] ^ IN[56] ^ IN[57] ^ IN[60] ^ IN[63] ^ IN[66] ^ IN[70] ^ IN[71] ^ IN[76] ^ IN[77] ^ IN[78] ^ IN[79] ^ IN[85] ^ IN[88] ^ IN[90] ^ IN[92] ^ IN[93] ^ IN[94] ^ IN[101] ^ IN[104] ^ IN[105] ^ IN[108] ^ IN[110] ^ IN[117] ^ IN[121] ^ IN[122] ^ IN[127] ^ IN[128] ^ IN[133] ^ IN[134] ^ IN[137] ^ IN[138] ^ IN[139] ^ IN[143] ^ IN[144] ^ IN[145] ^ IN[146] ^ IN[147] ^ IN[148] ^ IN[152] ^ IN[156] ^ IN[158] ^ IN[159] ^ IN[160] ^ IN[161] ^ IN[163] ^ IN[165] ^ IN[167] ^ IN[168] ^ IN[169] ^ IN[170] ^ IN[174] ^ IN[176] ^ IN[180] ^ IN[181] ^ IN[183] ^ IN[186] ^ IN[189] ^ IN[190] ^ IN[191] ^ IN[193] ^ IN[195] ^ IN[198] ^ IN[199] ^ IN[201] ^ IN[202] ^ IN[203] ^ IN[208] ^ IN[210] ^ IN[216] ^ IN[217] ^ IN[218] ^ IN[228] ^ IN[234] ^ IN[235] ^ IN[238] ^ IN[241] ^ IN[244] ^ IN[245] ^ IN[249] ^ IN[252] ^ IN[253] ^ IN[254] ^ CHK[2];
        SYN[3] = IN[0] ^ IN[2] ^ IN[4] ^ IN[6] ^ IN[9] ^ IN[10] ^ IN[11] ^ IN[13] ^ IN[14] ^ IN[15] ^ IN[16] ^ IN[19] ^ IN[21] ^ IN[25] ^ IN[26] ^ IN[28] ^ IN[29] ^ IN[32] ^ IN[34] ^ IN[35] ^ IN[37] ^ IN[42] ^ IN[45] ^ IN[46] ^ IN[47] ^ IN[48] ^ IN[49] ^ IN[55] ^ IN[56] ^ IN[63] ^ IN[69] ^ IN[71] ^ IN[78] ^ IN[80] ^ IN[81] ^ IN[82] ^ IN[83] ^ IN[85] ^ IN[86] ^ IN[87] ^ IN[88] ^ IN[95] ^ IN[96] ^ IN[99] ^ IN[102] ^ IN[108] ^ IN[110] ^ IN[111] ^ IN[113] ^ IN[114] ^ IN[115] ^ IN[116] ^ IN[117] ^ IN[118] ^ IN[123] ^ IN[131] ^ IN[133] ^ IN[134] ^ IN[143] ^ IN[146] ^ IN[152] ^ IN[153] ^ IN[154] ^ IN[155] ^ IN[156] ^ IN[157] ^ IN[158] ^ IN[160] ^ IN[161] ^ IN[163] ^ IN[164] ^ IN[166] ^ IN[168] ^ IN[170] ^ IN[172] ^ IN[173] ^ IN[175] ^ IN[178] ^ IN[179] ^ IN[180] ^ IN[182] ^ IN[183] ^ IN[186] ^ IN[190] ^ IN[194] ^ IN[195] ^ IN[201] ^ IN[206] ^ IN[210] ^ IN[213] ^ IN[222] ^ IN[226] ^ IN[227] ^ IN[229] ^ IN[230] ^ IN[231] ^ IN[232] ^ IN[240] ^ IN[241] ^ IN[242] ^ IN[248] ^ IN[249] ^ IN[251] ^ IN[252] ^ CHK[3];
        SYN[4] = IN[2] ^ IN[3] ^ IN[4] ^ IN[5] ^ IN[6] ^ IN[8] ^ IN[9] ^ IN[11] ^ IN[12] ^ IN[13] ^ IN[16] ^ IN[19] ^ IN[21] ^ IN[22] ^ IN[23] ^ IN[24] ^ IN[27] ^ IN[29] ^ IN[30] ^ IN[32] ^ IN[34] ^ IN[39] ^ IN[41] ^ IN[42] ^ IN[43] ^ IN[44] ^ IN[47] ^ IN[48] ^ IN[51] ^ IN[53] ^ IN[54] ^ IN[56] ^ IN[60] ^ IN[61] ^ IN[62] ^ IN[64] ^ IN[66] ^ IN[68] ^ IN[70] ^ IN[73] ^ IN[74] ^ IN[82] ^ IN[83] ^ IN[84] ^ IN[86] ^ IN[90] ^ IN[91] ^ IN[93] ^ IN[94] ^ IN[95] ^ IN[100] ^ IN[103] ^ IN[108] ^ IN[109] ^ IN[111] ^ IN[113] ^ IN[116] ^ IN[121] ^ IN[122] ^ IN[123] ^ IN[125] ^ IN[126] ^ IN[130] ^ IN[131] ^ IN[132] ^ IN[134] ^ IN[137] ^ IN[139] ^ IN[140] ^ IN[147] ^ IN[149] ^ IN[152] ^ IN[153] ^ IN[155] ^ IN[157] ^ IN[162] ^ IN[163] ^ IN[164] ^ IN[166] ^ IN[168] ^ IN[169] ^ IN[177] ^ IN[178] ^ IN[187] ^ IN[188] ^ IN[189] ^ IN[191] ^ IN[201] ^ IN[202] ^ IN[206] ^ IN[210] ^ IN[211] ^ IN[214] ^ IN[216] ^ IN[218] ^ IN[220] ^ IN[231] ^ IN[233] ^ IN[234] ^ IN[235] ^ IN[237] ^ IN[239] ^ IN[240] ^ IN[243] ^ IN[253] ^ CHK[4];
        SYN[5] = IN[2] ^ IN[3] ^ IN[7] ^ IN[8] ^ IN[13] ^ IN[14] ^ IN[15] ^ IN[17] ^ IN[20] ^ IN[24] ^ IN[25] ^ IN[27] ^ IN[28] ^ IN[30] ^ IN[31] ^ IN[35] ^ IN[36] ^ IN[37] ^ IN[38] ^ IN[39] ^ IN[40] ^ IN[47] ^ IN[52] ^ IN[53] ^ IN[55] ^ IN[56] ^ IN[57] ^ IN[61] ^ IN[63] ^ IN[69] ^ IN[71] ^ IN[74] ^ IN[75] ^ IN[77] ^ IN[79] ^ IN[88] ^ IN[89] ^ IN[90] ^ IN[95] ^ IN[98] ^ IN[99] ^ IN[100] ^ IN[103] ^ IN[106] ^ IN[107] ^ IN[113] ^ IN[118] ^ IN[119] ^ IN[124] ^ IN[126] ^ IN[127] ^ IN[128] ^ IN[130] ^ IN[131] ^ IN[139] ^ IN[140] ^ IN[141] ^ IN[147] ^ IN[148] ^ IN[150] ^ IN[151] ^ IN[153] ^ IN[154] ^ IN[158] ^ IN[159] ^ IN[161] ^ IN[162] ^ IN[163] ^ IN[166] ^ IN[168] ^ IN[170] ^ IN[172] ^ IN[175] ^ IN[176] ^ IN[183] ^ IN[184] ^ IN[186] ^ IN[189] ^ IN[191] ^ IN[195] ^ IN[205] ^ IN[207] ^ IN[213] ^ IN[215] ^ IN[217] ^ IN[218] ^ IN[221] ^ IN[224] ^ IN[225] ^ IN[226] ^ IN[228] ^ IN[230] ^ IN[234] ^ IN[238] ^ IN[243] ^ IN[244] ^ IN[245] ^ IN[246] ^ IN[247] ^ IN[248] ^ IN[249] ^ IN[251] ^ IN[255] ^ CHK[5];
        SYN[6] = IN[1] ^ IN[2] ^ IN[3] ^ IN[6] ^ IN[8] ^ IN[9] ^ IN[10] ^ IN[11] ^ IN[15] ^ IN[19] ^ IN[20] ^ IN[21] ^ IN[22] ^ IN[24] ^ IN[28] ^ IN[29] ^ IN[30] ^ IN[37] ^ IN[38] ^ IN[39] ^ IN[41] ^ IN[42] ^ IN[43] ^ IN[44] ^ IN[46] ^ IN[53] ^ IN[54] ^ IN[55] ^ IN[56] ^ IN[58] ^ IN[59] ^ IN[60] ^ IN[61] ^ IN[63] ^ IN[70] ^ IN[71] ^ IN[76] ^ IN[78] ^ IN[82] ^ IN[83] ^ IN[84] ^ IN[85] ^ IN[87] ^ IN[88] ^ IN[89] ^ IN[90] ^ IN[91] ^ IN[94] ^ IN[96] ^ IN[97] ^ IN[98] ^ IN[101] ^ IN[104] ^ IN[106] ^ IN[108] ^ IN[110] ^ IN[114] ^ IN[116] ^ IN[118] ^ IN[119] ^ IN[121] ^ IN[123] ^ IN[124] ^ IN[127] ^ IN[129] ^ IN[130] ^ IN[131] ^ IN[133] ^ IN[134] ^ IN[135] ^ IN[140] ^ IN[143] ^ IN[145] ^ IN[146] ^ IN[147] ^ IN[149] ^ IN[150] ^ IN[151] ^ IN[157] ^ IN[159] ^ IN[162] ^ IN[166] ^ IN[175] ^ IN[177] ^ IN[181] ^ IN[185] ^ IN[188] ^ IN[191] ^ IN[192] ^ IN[193] ^ IN[196] ^ IN[197] ^ IN[200] ^ IN[204] ^ IN[207] ^ IN[211] ^ IN[212] ^ IN[215] ^ IN[217] ^ IN[219] ^ IN[221] ^ IN[228] ^ IN[229] ^ IN[230] ^ IN[231] ^ IN[232] ^ IN[236] ^ IN[242] ^ IN[252] ^ CHK[6];
        SYN[7] = IN[2] ^ IN[5] ^ IN[6] ^ IN[7] ^ IN[8] ^ IN[10] ^ IN[12] ^ IN[14] ^ IN[15] ^ IN[18] ^ IN[19] ^ IN[22] ^ IN[23] ^ IN[24] ^ IN[26] ^ IN[27] ^ IN[28] ^ IN[31] ^ IN[34] ^ IN[35] ^ IN[37] ^ IN[38] ^ IN[44] ^ IN[46] ^ IN[47] ^ IN[48] ^ IN[53] ^ IN[58] ^ IN[59] ^ IN[64] ^ IN[65] ^ IN[67] ^ IN[70] ^ IN[72] ^ IN[74] ^ IN[75] ^ IN[76] ^ IN[77] ^ IN[78] ^ IN[79] ^ IN[82] ^ IN[83] ^ IN[88] ^ IN[90] ^ IN[91] ^ IN[92] ^ IN[93] ^ IN[94] ^ IN[96] ^ IN[97] ^ IN[99] ^ IN[101] ^ IN[103] ^ IN[105] ^ IN[106] ^ IN[107] ^ IN[108] ^ IN[110] ^ IN[111] ^ IN[112] ^ IN[115] ^ IN[117] ^ IN[119] ^ IN[120] ^ IN[122] ^ IN[124] ^ IN[126] ^ IN[128] ^ IN[129] ^ IN[134] ^ IN[136] ^ IN[139] ^ IN[141] ^ IN[144] ^ IN[145] ^ IN[150] ^ IN[151] ^ IN[154] ^ IN[161] ^ IN[162] ^ IN[164] ^ IN[165] ^ IN[167] ^ IN[170] ^ IN[171] ^ IN[173] ^ IN[181] ^ IN[185] ^ IN[187] ^ IN[188] ^ IN[190] ^ IN[193] ^ IN[194] ^ IN[196] ^ IN[206] ^ IN[209] ^ IN[210] ^ IN[212] ^ IN[213] ^ IN[215] ^ IN[218] ^ IN[219] ^ IN[224] ^ IN[226] ^ IN[229] ^ IN[231] ^ IN[233] ^ IN[234] ^ IN[235] ^ IN[238] ^ IN[240] ^ IN[243] ^ IN[246] ^ IN[247] ^ IN[248] ^ IN[255] ^ CHK[7];
        SYN[8] = IN[0] ^ IN[1] ^ IN[2] ^ IN[6] ^ IN[7] ^ IN[9] ^ IN[10] ^ IN[12] ^ IN[17] ^ IN[20] ^ IN[21] ^ IN[24] ^ IN[25] ^ IN[26] ^ IN[27] ^ IN[30] ^ IN[38] ^ IN[39] ^ IN[42] ^ IN[45] ^ IN[47] ^ IN[48] ^ IN[49] ^ IN[51] ^ IN[52] ^ IN[55] ^ IN[56] ^ IN[61] ^ IN[62] ^ IN[63] ^ IN[64] ^ IN[65] ^ IN[69] ^ IN[70] ^ IN[71] ^ IN[73] ^ IN[74] ^ IN[75] ^ IN[81] ^ IN[83] ^ IN[84] ^ IN[89] ^ IN[95] ^ IN[96] ^ IN[97] ^ IN[100] ^ IN[101] ^ IN[103] ^ IN[104] ^ IN[105] ^ IN[107] ^ IN[109] ^ IN[111] ^ IN[112] ^ IN[114] ^ IN[116] ^ IN[120] ^ IN[121] ^ IN[125] ^ IN[128] ^ IN[135] ^ IN[138] ^ IN[141] ^ IN[145] ^ IN[146] ^ IN[148] ^ IN[149] ^ IN[151] ^ IN[155] ^ IN[157] ^ IN[159] ^ IN[162] ^ IN[165] ^ IN[168] ^ IN[169] ^ IN[170] ^ IN[172] ^ IN[174] ^ IN[179] ^ IN[181] ^ IN[186] ^ IN[198] ^ IN[201] ^ IN[202] ^ IN[203] ^ IN[207] ^ IN[208] ^ IN[211] ^ IN[213] ^ IN[215] ^ IN[219] ^ IN[221] ^ IN[223] ^ IN[224] ^ IN[232] ^ IN[233] ^ IN[235] ^ IN[238] ^ IN[239] ^ IN[240] ^ IN[245] ^ IN[250] ^ CHK[8];
        SYN[9] = IN[0] ^ IN[1] ^ IN[3] ^ IN[8] ^ IN[9] ^ IN[13] ^ IN[15] ^ IN[17] ^ IN[19] ^ IN[23] ^ IN[24] ^ IN[26] ^ IN[28] ^ IN[30] ^ IN[31] ^ IN[32] ^ IN[33] ^ IN[34] ^ IN[39] ^ IN[41] ^ IN[42] ^ IN[44] ^ IN[45] ^ IN[48] ^ IN[49] ^ IN[51] ^ IN[53] ^ IN[54] ^ IN[58] ^ IN[60] ^ IN[61] ^ IN[62] ^ IN[65] ^ IN[66] ^ IN[67] ^ IN[69] ^ IN[71] ^ IN[74] ^ IN[78] ^ IN[79] ^ IN[81] ^ IN[82] ^ IN[83] ^ IN[91] ^ IN[92] ^ IN[98] ^ IN[99] ^ IN[101] ^ IN[103] ^ IN[106] ^ IN[107] ^ IN[112] ^ IN[115] ^ IN[116] ^ IN[118] ^ IN[121] ^ IN[125] ^ IN[128] ^ IN[133] ^ IN[136] ^ IN[139] ^ IN[142] ^ IN[143] ^ IN[144] ^ IN[149] ^ IN[150] ^ IN[154] ^ IN[155] ^ IN[157] ^ IN[159] ^ IN[160] ^ IN[161] ^ IN[163] ^ IN[173] ^ IN[178] ^ IN[180] ^ IN[182] ^ IN[187] ^ IN[189] ^ IN[193] ^ IN[195] ^ IN[197] ^ IN[198] ^ IN[200] ^ IN[205] ^ IN[207] ^ IN[209] ^ IN[210] ^ IN[212] ^ IN[214] ^ IN[215] ^ IN[216] ^ IN[225] ^ IN[226] ^ IN[227] ^ IN[228] ^ IN[229] ^ IN[233] ^ IN[237] ^ IN[238] ^ IN[239] ^ IN[249] ^ IN[250] ^ IN[254] ^ CHK[9];
        SYN[10] = IN[0] ^ IN[1] ^ IN[2] ^ IN[5] ^ IN[6] ^ IN[8] ^ IN[9] ^ IN[10] ^ IN[11] ^ IN[12] ^ IN[14] ^ IN[16] ^ IN[17] ^ IN[19] ^ IN[22] ^ IN[23] ^ IN[24] ^ IN[25] ^ IN[27] ^ IN[28] ^ IN[29] ^ IN[31] ^ IN[33] ^ IN[34] ^ IN[35] ^ IN[36] ^ IN[45] ^ IN[46] ^ IN[47] ^ IN[49] ^ IN[50] ^ IN[51] ^ IN[55] ^ IN[57] ^ IN[58] ^ IN[59] ^ IN[60] ^ IN[62] ^ IN[65] ^ IN[67] ^ IN[68] ^ IN[70] ^ IN[71] ^ IN[72] ^ IN[78] ^ IN[82] ^ IN[83] ^ IN[84] ^ IN[86] ^ IN[87] ^ IN[92] ^ IN[93] ^ IN[94] ^ IN[99] ^ IN[100] ^ IN[103] ^ IN[105] ^ IN[106] ^ IN[107] ^ IN[108] ^ IN[110] ^ IN[112] ^ IN[116] ^ IN[117] ^ IN[118] ^ IN[119] ^ IN[120] ^ IN[127] ^ IN[129] ^ IN[130] ^ IN[132] ^ IN[133] ^ IN[142] ^ IN[143] ^ IN[145] ^ IN[146] ^ IN[155] ^ IN[157] ^ IN[164] ^ IN[166] ^ IN[169] ^ IN[174] ^ IN[176] ^ IN[177] ^ IN[180] ^ IN[182] ^ IN[183] ^ IN[184] ^ IN[189] ^ IN[193] ^ IN[194] ^ IN[197] ^ IN[200] ^ IN[204] ^ IN[205] ^ IN[206] ^ IN[207] ^ IN[220] ^ IN[222] ^ IN[224] ^ IN[228] ^ IN[229] ^ IN[237] ^ IN[245] ^ IN[250] ^ IN[251] ^ IN[255] ^ CHK[10];
        SYN[11] = IN[0] ^ IN[4] ^ IN[6] ^ IN[10] ^ IN[11] ^ IN[15] ^ IN[17] ^ IN[19] ^ IN[21] ^ IN[22] ^ IN[26] ^ IN[27] ^ IN[28] ^ IN[30] ^ IN[31] ^ IN[32] ^ IN[34] ^ IN[35] ^ IN[36] ^ IN[37] ^ IN[40] ^ IN[41] ^ IN[43] ^ IN[44] ^ IN[45] ^ IN[50] ^ IN[51] ^ IN[52] ^ IN[53] ^ IN[54] ^ IN[56] ^ IN[57] ^ IN[58] ^ IN[65] ^ IN[67] ^ IN[73] ^ IN[75] ^ IN[76] ^ IN[77] ^ IN[78] ^ IN[79] ^ IN[80] ^ IN[84] ^ IN[87] ^ IN[90] ^ IN[92] ^ IN[94] ^ IN[98] ^ IN[99] ^ IN[101] ^ IN[105] ^ IN[106] ^ IN[108] ^ IN[111] ^ IN[113] ^ IN[114] ^ IN[115] ^ IN[117] ^ IN[122] ^ IN[126] ^ IN[128] ^ IN[129] ^ IN[132] ^ IN[135] ^ IN[140] ^ IN[143] ^ IN[151] ^ IN[152] ^ IN[155] ^ IN[157] ^ IN[158] ^ IN[161] ^ IN[163] ^ IN[167] ^ IN[170] ^ IN[171] ^ IN[172] ^ IN[173] ^ IN[179] ^ IN[180] ^ IN[182] ^ IN[183] ^ IN[192] ^ IN[193] ^ IN[199] ^ IN[202] ^ IN[203] ^ IN[204] ^ IN[206] ^ IN[208] ^ IN[209] ^ IN[210] ^ IN[212] ^ IN[213] ^ IN[214] ^ IN[215] ^ IN[216] ^ IN[219] ^ IN[221] ^ IN[227] ^ IN[231] ^ IN[233] ^ IN[241] ^ IN[242] ^ IN[247] ^ IN[250] ^ IN[254] ^ IN[255] ^ CHK[11];
        SYN[12] = IN[2] ^ IN[3] ^ IN[4] ^ IN[9] ^ IN[11] ^ IN[12] ^ IN[15] ^ IN[18] ^ IN[19] ^ IN[20] ^ IN[23] ^ IN[28] ^ IN[29] ^ IN[32] ^ IN[35] ^ IN[39] ^ IN[40] ^ IN[43] ^ IN[45] ^ IN[46] ^ IN[48] ^ IN[50] ^ IN[52] ^ IN[53] ^ IN[54] ^ IN[56] ^ IN[58] ^ IN[61] ^ IN[62] ^ IN[63] ^ IN[65] ^ IN[66] ^ IN[69] ^ IN[70] ^ IN[73] ^ IN[75] ^ IN[76] ^ IN[77] ^ IN[81] ^ IN[82] ^ IN[84] ^ IN[85] ^ IN[86] ^ IN[90] ^ IN[93] ^ IN[95] ^ IN[96] ^ IN[97] ^ IN[98] ^ IN[101] ^ IN[102] ^ IN[103] ^ IN[104] ^ IN[108] ^ IN[109] ^ IN[111] ^ IN[116] ^ IN[119] ^ IN[120] ^ IN[122] ^ IN[127] ^ IN[131] ^ IN[132] ^ IN[135] ^ IN[137] ^ IN[138] ^ IN[139] ^ IN[142] ^ IN[143] ^ IN[149] ^ IN[150] ^ IN[156] ^ IN[158] ^ IN[160] ^ IN[161] ^ IN[165] ^ IN[168] ^ IN[169] ^ IN[170] ^ IN[171] ^ IN[173] ^ IN[176] ^ IN[179] ^ IN[182] ^ IN[183] ^ IN[184] ^ IN[188] ^ IN[189] ^ IN[192] ^ IN[195] ^ IN[196] ^ IN[199] ^ IN[200] ^ IN[206] ^ IN[208] ^ IN[212] ^ IN[214] ^ IN[217] ^ IN[221] ^ IN[222] ^ IN[225] ^ IN[230] ^ IN[231] ^ IN[232] ^ IN[233] ^ IN[236] ^ IN[240] ^ IN[242] ^ IN[243] ^ IN[248] ^ IN[255] ^ CHK[12];
        SYN[13] = IN[1] ^ IN[3] ^ IN[4] ^ IN[5] ^ IN[6] ^ IN[7] ^ IN[13] ^ IN[14] ^ IN[17] ^ IN[18] ^ IN[20] ^ IN[23] ^ IN[24] ^ IN[29] ^ IN[30] ^ IN[31] ^ IN[33] ^ IN[35] ^ IN[39] ^ IN[40] ^ IN[41] ^ IN[45] ^ IN[49] ^ IN[50] ^ IN[52] ^ IN[53] ^ IN[55] ^ IN[58] ^ IN[59] ^ IN[61] ^ IN[64] ^ IN[67] ^ IN[68] ^ IN[69] ^ IN[71] ^ IN[72] ^ IN[75] ^ IN[76] ^ IN[80] ^ IN[82] ^ IN[83] ^ IN[85] ^ IN[86] ^ IN[88] ^ IN[89] ^ IN[91] ^ IN[94] ^ IN[95] ^ IN[97] ^ IN[98] ^ IN[107] ^ IN[109] ^ IN[110] ^ IN[112] ^ IN[114] ^ IN[115] ^ IN[119] ^ IN[120] ^ IN[121] ^ IN[122] ^ IN[123] ^ IN[126] ^ IN[131] ^ IN[135] ^ IN[141] ^ IN[142] ^ IN[143] ^ IN[145] ^ IN[150] ^ IN[151] ^ IN[152] ^ IN[154] ^ IN[155] ^ IN[158] ^ IN[165] ^ IN[172] ^ IN[174] ^ IN[175] ^ IN[177] ^ IN[182] ^ IN[185] ^ IN[187] ^ IN[192] ^ IN[195] ^ IN[196] ^ IN[198] ^ IN[199] ^ IN[204] ^ IN[207] ^ IN[209] ^ IN[214] ^ IN[222] ^ IN[223] ^ IN[232] ^ IN[234] ^ IN[237] ^ IN[239] ^ IN[244] ^ IN[247] ^ IN[251] ^ IN[254] ^ CHK[13];
        SYN[14] = IN[0] ^ IN[1] ^ IN[2] ^ IN[4] ^ IN[12] ^ IN[15] ^ IN[20] ^ IN[25] ^ IN[29] ^ IN[32] ^ IN[33] ^ IN[35] ^ IN[37] ^ IN[38] ^ IN[41] ^ IN[43] ^ IN[44] ^ IN[48] ^ IN[50] ^ IN[51] ^ IN[53] ^ IN[55] ^ IN[56] ^ IN[59] ^ IN[61] ^ IN[64] ^ IN[67] ^ IN[68] ^ IN[69] ^ IN[73] ^ IN[77] ^ IN[79] ^ IN[83] ^ IN[84] ^ IN[87] ^ IN[88] ^ IN[91] ^ IN[93] ^ IN[94] ^ IN[98] ^ IN[100] ^ IN[102] ^ IN[103] ^ IN[104] ^ IN[105] ^ IN[106] ^ IN[111] ^ IN[114] ^ IN[115] ^ IN[116] ^ IN[117] ^ IN[118] ^ IN[125] ^ IN[126] ^ IN[129] ^ IN[130] ^ IN[133] ^ IN[141] ^ IN[144] ^ IN[145] ^ IN[148] ^ IN[151] ^ IN[153] ^ IN[155] ^ IN[159] ^ IN[160] ^ IN[161] ^ IN[162] ^ IN[163] ^ IN[164] ^ IN[165] ^ IN[171] ^ IN[172] ^ IN[176] ^ IN[178] ^ IN[180] ^ IN[182] ^ IN[186] ^ IN[189] ^ IN[190] ^ IN[191] ^ IN[192] ^ IN[193] ^ IN[196] ^ IN[197] ^ IN[198] ^ IN[201] ^ IN[206] ^ IN[207] ^ IN[208] ^ IN[211] ^ IN[212] ^ IN[213] ^ IN[217] ^ IN[219] ^ IN[223] ^ IN[225] ^ IN[226] ^ IN[227] ^ IN[230] ^ IN[231] ^ IN[233] ^ IN[234] ^ IN[246] ^ IN[251] ^ IN[252] ^ IN[253] ^ CHK[14];
        SYN[15] = IN[1] ^ IN[7] ^ IN[11] ^ IN[12] ^ IN[13] ^ IN[15] ^ IN[18] ^ IN[20] ^ IN[23] ^ IN[24] ^ IN[25] ^ IN[26] ^ IN[32] ^ IN[35] ^ IN[36] ^ IN[38] ^ IN[39] ^ IN[40] ^ IN[42] ^ IN[44] ^ IN[47] ^ IN[48] ^ IN[50] ^ IN[51] ^ IN[52] ^ IN[54] ^ IN[58] ^ IN[62] ^ IN[67] ^ IN[68] ^ IN[70] ^ IN[71] ^ IN[72] ^ IN[74] ^ IN[76] ^ IN[78] ^ IN[79] ^ IN[80] ^ IN[82] ^ IN[85] ^ IN[86] ^ IN[88] ^ IN[91] ^ IN[92] ^ IN[97] ^ IN[99] ^ IN[101] ^ IN[102] ^ IN[104] ^ IN[105] ^ IN[110] ^ IN[111] ^ IN[112] ^ IN[113] ^ IN[118] ^ IN[128] ^ IN[129] ^ IN[130] ^ IN[131] ^ IN[136] ^ IN[137] ^ IN[138] ^ IN[142] ^ IN[143] ^ IN[147] ^ IN[148] ^ IN[150] ^ IN[151] ^ IN[155] ^ IN[164] ^ IN[165] ^ IN[168] ^ IN[178] ^ IN[180] ^ IN[183] ^ IN[184] ^ IN[185] ^ IN[188] ^ IN[190] ^ IN[192] ^ IN[203] ^ IN[210] ^ IN[213] ^ IN[215] ^ IN[217] ^ IN[218] ^ IN[220] ^ IN[223] ^ IN[224] ^ IN[231] ^ IN[236] ^ IN[239] ^ IN[241] ^ IN[246] ^ IN[247] ^ IN[250] ^ IN[253] ^ IN[254] ^ CHK[15];

       ERR = |SYN;
       SGL = ^SYN & ERR;
       DBL = ~^SYN & ERR;
    end

corrector corr_mod (.IN(IN), .SYN(SYN), .OUT(OUT));

endmodule



